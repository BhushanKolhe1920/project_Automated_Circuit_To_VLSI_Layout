MACRO AND4
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND4 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal1 ;
        RECT 0.00000000 30500.00000000 48000.00000000 33500.00000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal1 ;
        RECT 0.00000000 -1500.00000000 48000.00000000 1500.00000000 ;
    END
  END GND

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 7000.00000000 9500.00000000 9000.00000000 11500.00000000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 15000.00000000 9500.00000000 17000.00000000 11500.00000000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 23000.00000000 9500.00000000 25000.00000000 11500.00000000 ;
    END
  END C

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 31000.00000000 9500.00000000 33000.00000000 11500.00000000 ;
    END
  END D

  PIN Z
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 43000.00000000 8500.00000000 45000.00000000 10500.00000000 ;
    END
  END Z


END AND4
